
module RefModule (
  input a,
  input b,
  input c,
  input d,
  output dout,
  output out_n
);

  wire w1, w2;
  assign w1 = a&b;
  assign w2 = c&d;
  assign dout = w1|w2;
  assign out_n = ~dout;

endmodule

