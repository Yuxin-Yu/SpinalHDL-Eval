
module RefModule (
  input din,
  output dout
);

  assign dout = din;

endmodule

