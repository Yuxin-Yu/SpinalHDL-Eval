
module RefModule (
  output dout
);

  assign dout = 1'b0;

endmodule

